
`include "common.v"

module control (
    input                   	    instr_valid,
    input [`INSTR_WIDTH - 1: 0]     instr,

    output 	reg	[`BRANCH_TYPE_BUS]  branch,
    output  reg	            	    mem_read,
    output  reg	            	    mem2reg,
    output  reg	            	    mem_write,
    output  reg	            	    reg_write,
    output  reg	                    unknown_op,
    output  reg	            	    ALU_in1_type,
    output  reg	[`ALU_IN2_BUS] 	    ALU_in2_type,
    output  reg	[`ALUOP_BUS]	    ALU_OP,
    output  reg [`INSTR_TYPE_BUS]   instr_type,
    output  reg                     stall,                        
    output  reg [`OP_WIDTH_BUS]     op_width
);

    always @(*) begin
        if (instr_valid == `FALSE)                                  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_NULL; instr_type = `NULL_TYPE;	op_width = `OP_WIDTH_8_REG; stall = `FALSE; unknown_op = `FALSE;    end
        else begin
            casez (instr)                                           
                32'bzzzzzzzzzzzz_zzzzz_000_zzzzz__0010011/*addi */: begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;				            end
                32'bzzzzzzzzzzzzzzzzzzzz_zzzzz____0010111/*auipc*/: begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_PC;  ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `U_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;          				end
                32'bzzzzzzzzzzzzzzzzzzzz_zzzzz____1101111/*jal*/:   begin branch = `BRANCH_JAL;  mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_PC;  ALU_in2_type = `ALU_IN2_4;    ALU_OP = `ALUOP_ADD;  instr_type = `J_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;           				end
                32'bzzzzzzz_zzzzz_zzzzz_011_zzzzz_0100011/*sd*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_1; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `S_TYPE;   	op_width = `OP_WIDTH_8_MEM; stall = `TRUE;		    				end
                32'bzzzzzzzzzzzz_zzzzz_000_zzzzz__1100111/*jalr*/:  begin branch = `BRANCH_JALR; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_PC;  ALU_in2_type = `ALU_IN2_4;    ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;           				end
                32'bzzzzzzzzzzzz_zzzzz_011_zzzzz__0000011/*ld*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_1; mem2reg = `ENA_1; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;   	op_width = `OP_WIDTH_8_MEM; stall = `TRUE;							end
                32'b0000000_zzzzz_zzzzz_000_zzzzz_0110011/*add*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_ADD;  instr_type = `R_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;          				end
                32'b0100000_zzzzz_zzzzz_000_zzzzz_0110011/*sub*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SUB;  instr_type = `R_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;           				end
                32'bzzzzzzzzzzzz_zzzzz_011_zzzzz__0010011/*sltiu*/: begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_UL;   instr_type = `I_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;           				end
                32'bzzzzzzz_zzzzz_zzzzz_000_zzzzz_1100011/*beq*/:   begin branch = `BRANCH_BEQ;  mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SUB;  instr_type = `B_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;           				end
                32'bzzzzzzz_zzzzz_zzzzz_001_zzzzz_1100011/*bne*/:   begin branch = `BRANCH_BNE;  mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SUB;  instr_type = `B_TYPE;   	op_width = `OP_WIDTH_8_REG; stall = `FALSE;           				end
                32'bzzzzzzzzzzzz_zzzzz_000_zzzzz__0011011/*addiw*/: begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;         				end
                32'bzzzzzzzzzzzz_zzzzz_010_zzzzz__0000011/*lw*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_1; mem2reg = `ENA_1; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;   	op_width = `OP_WIDTH_4_MEM; stall = `TRUE;                          end
                32'b0000000_zzzzz_zzzzz_000_zzzzz_0111011/*addw*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_ADD;  instr_type = `R_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;        				    end
                32'bzzzzzzz_zzzzz_zzzzz_001_zzzzz_0100011/*sh*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_1; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `S_TYPE;    op_width = `OP_WIDTH_2_MEM; stall = `TRUE;        				    end
                32'b010000_zzzzzz_zzzzz_101_zzzzz_0010011/*srai*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_SRAI; instr_type = `I_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzzzzzzz_zzzzz_100_zzzzz__0000011/*lbu*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_1; mem2reg = `ENA_1; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_1_MEM; stall = `TRUE;        				    end
                32'bzzzzzzzzzzzz_zzzzz_111_zzzzz__0010011/*andi*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_AND;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b0000000_zzzzz_zzzzz_001_zzzzz_0111011/*sllw*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SLLW; instr_type = `R_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;        				    end
                32'b0000000_zzzzz_zzzzz_111_zzzzz_0110011/*and*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_AND;  instr_type = `R_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b0000000_zzzzz_zzzzz_011_zzzzz_0110011/*sltu*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_UL;   instr_type = `R_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzzzzzzz_zzzzz_100_zzzzz__0010011/*xori*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_XOR;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b0000000_zzzzz_zzzzz_110_zzzzz_0110011/*or*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_OR;   instr_type = `R_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzz_zzzzz_zzzzz_000_zzzzz_0100011/*sb*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_1; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `S_TYPE;    op_width = `OP_WIDTH_1_MEM; stall = `TRUE;        				    end
                32'b000000_zzzzzz_zzzzz_001_zzzzz_0010011/*slli*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_SLLI; instr_type = `I_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b000000_zzzzzz_zzzzz_101_zzzzz_0010011/*srli*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_SRL;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzz_zzzzz_zzzzz_101_zzzzz_1100011/*bge*/:   begin branch = `BRANCH_BGE;  mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SUB;  instr_type = `B_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzz_zzzzz_zzzzz_010_zzzzz_0100011/*sw*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_1; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `S_TYPE;    op_width = `OP_WIDTH_4_MEM; stall = `TRUE;        				    end
                32'bzzzzzzz_zzzzz_zzzzz_100_zzzzz_1100011/*blt*/:   begin branch = `BRANCH_BLT;  mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SUB;  instr_type = `B_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzz_zzzzz_zzzzz_111_zzzzz_1100011/*bgeu*/:  begin branch = `BRANCH_BGEU; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_GEU;  instr_type = `B_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzz_zzzzz_zzzzz_110_zzzzz_1100011/*bltu*/:  begin branch = `BRANCH_BLTU; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_LTU;  instr_type = `B_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b000000_zzzzz_zzzzz_010_zzzzz__0110011/*slt*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SLT;  instr_type = `R_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzzzzzzz_zzzzz_001_zzzzz__0000011/*lh*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_1; mem2reg = `ENA_1; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_2_MEM; stall = `TRUE;        				    end
                32'bzzzzzzzzzzzz_zzzzz_101_zzzzz__0000011/*lhu*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_1; mem2reg = `ENA_1; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_2_MEM; stall = `TRUE;        				    end
                32'b0100000_zzzzz_zzzzz_000_zzzzz_0111011/*subw*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SUB;  instr_type = `R_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;        				    end
                32'b000000_zzzzzz_zzzzz_001_zzzzz_0011011/*slliw*/: begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_SLLI; instr_type = `I_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;        				    end
                32'b010000_zzzzzz_zzzzz_101_zzzzz_0011011/*sraiw*/: begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_SRAW; instr_type = `I_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;        				    end
                32'bzzzzzzzzzzzzzzzzzzzz_zzzzz____0110111/*lui*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_MV2;  instr_type = `U_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b000000_zzzzzz_zzzzz_101_zzzzz_0011011/*srliw*/: begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_SRLIW;instr_type = `I_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;        				    end
                32'b0100000_zzzzz_zzzzz_101_zzzzz_0111011/*sraw*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SRAW; instr_type = `R_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;        				    end
                32'b0000000_zzzzz_zzzzz_101_zzzzz_0111011/*srlw*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SRLW; instr_type = `R_TYPE;    op_width = `OP_WIDTH_4_REG; stall = `FALSE;        				    end
                32'bzzzzzzz_zzzzz_zzzzz_110_zzzzz_0010011/*ori*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_OR;   instr_type = `I_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzzzzzzz_zzzzz_000_zzzzz__0000011/*lb*/:    begin branch = `BRANCH_NULL; mem_read = `ENA_1; mem2reg = `ENA_1; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_1_MEM; stall = `TRUE;        				    end
                32'bzzzzzzzzzzzz_zzzzz_110_zzzzz__0000011/*lwu*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_1; mem2reg = `ENA_1; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_ADD;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_4_MEM; stall = `TRUE;        				    end
                32'b0000000_zzzzz_zzzzz_001_zzzzz_0110011/*sll*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SLL;  instr_type = `R_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'bzzzzzzzzzzzz_zzzzz_010_zzzzz__0010011/*slti*/:  begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_SIMM; ALU_OP = `ALUOP_SLT;  instr_type = `I_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b0100000_zzzzz_zzzzz_101_zzzzz_0110011/*sra*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SRA;  instr_type = `R_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b0000000_zzzzz_zzzzz_101_zzzzz_0110011/*srl*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_SRL;  instr_type = `R_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                32'b0000000_zzzzz_zzzzz_100_zzzzz_0110011/*xor*/:   begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_1; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_XOR;  instr_type = `R_TYPE;    op_width = `OP_WIDTH_8_REG; stall = `FALSE;        				    end
                default:                                            begin branch = `BRANCH_NULL; mem_read = `ENA_0; mem2reg = `ENA_0; mem_write = `ENA_0; reg_write = `ENA_0; ALU_in1_type = `ALU_IN1_REG; ALU_in2_type = `ALU_IN2_REG;  ALU_OP = `ALUOP_NULL; instr_type = `NULL_TYPE; op_width = `OP_WIDTH_8_REG;                 unknown_op = `TRUE;     end
            endcase
        end
    end

endmodule
